// если нажата кнопка, то горит светодиод 4
module top(
    input A,
    output LED4
);
assign LED4 = A;
endmodule
