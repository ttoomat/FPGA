module gw_gao(
    clk,
    \t1/data_ind[2] ,
    \t1/data_ind[1] ,
    \t1/data_ind[0] ,
    \t1/tx ,
    \t1/trig ,
    \t1/present_state[1] ,
    \t1/present_state[0] ,
    \t1/next_state[1] ,
    \t1/next_state[0] ,
    \data1[7] ,
    \data1[6] ,
    \data1[5] ,
    \data1[4] ,
    \data1[3] ,
    \data1[2] ,
    \data1[1] ,
    \data1[0] ,
    \t1/reset ,
    \t1/tc ,
    iclk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input clk;
input \t1/data_ind[2] ;
input \t1/data_ind[1] ;
input \t1/data_ind[0] ;
input \t1/tx ;
input \t1/trig ;
input \t1/present_state[1] ;
input \t1/present_state[0] ;
input \t1/next_state[1] ;
input \t1/next_state[0] ;
input \data1[7] ;
input \data1[6] ;
input \data1[5] ;
input \data1[4] ;
input \data1[3] ;
input \data1[2] ;
input \data1[1] ;
input \data1[0] ;
input \t1/reset ;
input \t1/tc ;
input iclk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire clk;
wire \t1/data_ind[2] ;
wire \t1/data_ind[1] ;
wire \t1/data_ind[0] ;
wire \t1/tx ;
wire \t1/trig ;
wire \t1/present_state[1] ;
wire \t1/present_state[0] ;
wire \t1/next_state[1] ;
wire \t1/next_state[0] ;
wire \data1[7] ;
wire \data1[6] ;
wire \data1[5] ;
wire \data1[4] ;
wire \data1[3] ;
wire \data1[2] ;
wire \data1[1] ;
wire \data1[0] ;
wire \t1/reset ;
wire \t1/tc ;
wire iclk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top u_ao_top(
    .control(control0[9:0]),
    .data_i({clk,\t1/data_ind[2] ,\t1/data_ind[1] ,\t1/data_ind[0] ,\t1/tx ,\t1/trig ,\t1/present_state[1] ,\t1/present_state[0] ,\t1/next_state[1] ,\t1/next_state[0] ,\data1[7] ,\data1[6] ,\data1[5] ,\data1[4] ,\data1[3] ,\data1[2] ,\data1[1] ,\data1[0] ,\t1/reset ,\t1/tc }),
    .clk_i(iclk)
);

endmodule
