module top(
    input Power,
    output LED4
);
assign LED4 = Power;
endmodule
