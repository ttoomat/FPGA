module lut_top (
    input reg clk,

    input reg enable,
    input  reg S, A, B, C,
    output reg Z
);
/*
Сначала создайте 8-битный регистр сдвига с 8 D-триггерами.
Обозначьте выходы триггеров Q[0]...Q[7].
Вход регистра сдвига должен быть обозначен как S, он поступает на вход Q[0] (старший бит сдвигается первым).
Enable разрешает считать S.
Затем добавьте в схему 3 дополнительных входа A, B, C и выход Z.
Схема должна вести себя следующим образом: когда ABC равен 000, Z=Q[0], 
когда ABC равен 001, Z=Q[1] и так далее. 
Ваша схема должна содержать ТОЛЬКО 8-битный регистр сдвига и мультиплексоры.

Кроме создания LUT вам нужно определить 3 функции из testbench.
*/
reg out0;
// ниже - 8-битный регистр выходов с триггеров
reg [7:0]Q;
// должно быть: всё это запускается при изменении s

always @(posedge clk) begin
    // если enable - каждый такт сдвигаем S
    if (enable) begin
    Q[0] <= S;
    Q[1] <= Q[0];
    Q[2] <= Q[1];
    Q[3] <= Q[2];
    Q[4] <= Q[3];
    Q[5] <= Q[4];
    Q[6] <= Q[5];
    Q[7] <= Q[6];
    end
end

always @(*) begin
    case ({A, B, C})
    3'b000: Z = Q[0];
    3'b001: Z = Q[1];
    3'b010: Z = Q[2];
    3'b011: Z = Q[3];
    3'b100: Z = Q[4];
    3'b101: Z = Q[5];
    3'b110: Z = Q[6];
    3'b111: Z = Q[7];
    endcase
end

endmodule

/*
в каком смысле определить функции?
*/